-- Elementos de Sistemas
-- by Luciano Soares
-- Ram4K.vhd

Library ieee; 
use ieee.std_logic_1164.all;

  
entity Ram4K is
	port(
		clock   in  STD_LOGIC;
		input   in  STD_LOGIC_VECTOR(15 downto 0);
		load    in  STD_LOGIC;
		address in  STD_LOGIC_VECTOR(11 downto 0);
		output  out STD_LOGIC_VECTOR(15 downto 0)
	);
end entity;
